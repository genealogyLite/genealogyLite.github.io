10002||10001|Elizabeta I.|Kurjaković|Zrinski||||||||||
10004||10005|Ana I.|Zrinski|||1410||||||||
10006||10005|Margareta I.|Zrinski|||||||||||
10008|||Sofija|Zrinski|||||||||||
10010|||Jelena|Zrinski|Babonić||||||||princess of Blagaj||
10012||10007|Katarina I.|Zrinski|||||||||||
10014||10007|Klara|Zrinski|||||||||||
10016||10007|Margareta II.|Zrinski||3|1442|||1488|||||
10018||10007|Ilka|Zrinski||3|1442|||1488|||||
10030|10008|10019|Jelena|Karlović|Zrinski||||||||||
10032|10008|10019|Margareta|Zrinski|||||||||||
10034|||Jelena|Zrinski|Karlović||||||||||
10036|10034|10035|Jelena|Tahy|Zrinski||||||||||
10038|10034|10035|Margareta III.|Zrinski|||||||||||
10040|10034|10035|Katarina  |Zrinski|Fraknopan of Ozalj|||||1561|||||
10042|10034|10035|Eva|Zrinski|Rožemberk/Rosenberg||1537|||1501|||||
10050|10040|10045|Jelena|Zrinski|||1546|||1585|||||
10052|10040|10045|Katarina II.|Zrinski|||1548|||1585|||||
10054|10040|10045|Ana|Zrinski|d’Arco|||||1570|||||
10056|10040|10045|Sofija|Zrinski|Stubenberg||||||||||
10058|10040|10045|Doroteja|Zrinski|||1550|||1617|||||
10060|10040|10045|Uršula|Zrinski|||1552|||1593|||||
10062|10040|10045|Barbara|Zrinski|||1554||||||||
10064|10040|10045|Margareta IV.|Zrinski|||1555|||1588|||||
10066|10040|10045|Ana II.|Zrinski|||1557||||||||
10068|10040|10045|Magdalena|Zrinski|||1561||||||||
10070|10056|10053|Barbara|Zrinski|||||||||||
10072|10056|10053|Elizabeta II.|Erdődy|Zrinski||||||||||
10074|10056|10053|Suzana|Lenković|Zrinski||||||||||
10076|||Magdalena|Zrinski|Széchy||||||||||
10080|||Marija Euzebija|Zrinski|Drašković|||||1650|||||
10082|||Marija Sofija|Zrinski|Löbl|||||1676|||||
10084|||Ana Katarina|Zrinski|Frankopan of Tržac||1625||Bosiljevo|1673||Graz|||
10090|10082|10081|Marija Terezija Barbara|Zrinski|||1655|||1658|||||
10092|10082|10081|Marija Katarina|Zrinski|||1656||||||||
10094|||Marija Katarina |Zrinski|Lamberg||||||||||
10096|10084|10083|Jelena|Rákóczi|Zrinski||1643||Ozalj|1703||Nicomedia|||
10098|10084|10083|Judita Pertonila|Zrinski|||1652||Ozalj|1600||Zagreb|||
10100|10084|10083|Zora Veronika|Zrinski|||1658||Ozalj|1735||Klanenfurt|||
