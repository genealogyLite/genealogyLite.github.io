10002|10003||||||||
10010|10019||||||||
10008|10019||||||||
10030|10039||||||||
10034|10035||||||||
10036|10041||||||||
10038|10063||||||||
10040|10045||||||||
10042|10045||||||||
10054|10053||||||||
10056|10053||||||||
10072|10073||||||||
10074|10075||||||||
10076|10077||||||||
10080|10081||||||||
10082|10081||||||||
10084|10083||||||||
10094|10093||||||||
