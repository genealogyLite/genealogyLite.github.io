10001|||Juraj I.|Zrinski|1|1300|||1361||||House of Zrinski primogenitor|<zrinski.html#10001>
10003|||Toma|Kurjaković|3|1320|||1380|||||
10005||10001|Pavao I.|Zrinski||1357|||1414||Zagreb|||
10007||10005|Petar I.|Zrinski||1408|||1446|||||
10009||10005|Nikola I.|Zrinski|1|1400|||1439|||||
10015||10007|Mirko|Zrinski||1423|||1435|||||
10017||10007|Pavao II.|Zrinski||1429|||1449|||||
10019||10007|Petar II.|Zrinski||1435|||1493|252|Krbava Field||Died in the battle of Krbava|
10021||10007|Juraj II.|Zrinski||1435|||1480|||||
10023||10007|Martin|Zrinski||||||||||
10031|10008|10019|Pavao III.|Zrinski||1465|||1493|252|Krbava Field||Died in the battle of Krbava|
10033|10008|10019|Bernard|Zrinski||||||||||
10035|10010|10019|Nikola III.|Zrinski||1489|||1534||Zrin|||
10037||10021|Nikola II.|Zrinski||||||||||
10041|||Ferenc|Tahy||||||||||
10049|10034|10035|Ivan I.|Zrinski||||||||||
10045|10034|10035|Nikola IV.|Zrinski|1|1508||Zrin|1566|250|Szigetvár|Ban of Croatia|Died in the siege of Szigetvár|<https://en.wikipedia.org/wiki/Nikola_IV_Zrinski>
10047|10034|10035|Petar III.|Zrinski||||||||||
10063|||Ivan|Alapić||||||||||
10043|10034|10035|Juraj III.|Zrinski||||||||||
10051|10040|10045|Ivan II.|Zrinski||||||||||
10053|10040|10045|Juraj IV.|Zrinski||||||||||
10055|10040|10045|Krsto|Zrinski||||||||||
10057|10040|10045|Vuk|Zrinski||||||||||
10059|10040|10045|Nikola V.|Zrinski||||||||||
10061|10042|10047|Ivan III.|Zrinski||||||||||
10071|10054|10053|Nikola VI |Zrinski||||||||||
10077|10056|10053|Juraj V.|Zrinski||||||||Ban of Croatia||
10073|||Toma|Erdödy||||||||||
10075|||Juraj|Lenković||||||||||
10081|10076|10077|Nikola VII.|Zrinski||||||||||
10083|10076|10077|Petar IV.|Zrinski||1621|157|Vrbovec|1671|120|Wiener Neustadt|Ban of Croatia|Executed by Habsburg monarchy |<https://en.wikipedia.org/wiki/Petar_Zrinski>
10091|10082|10081|Izak|Zrinski||||||||||
10093|10082|10081|Adam|Zrinski||||||||||
10095|10084|10083|Ivan IV. Antun|Zrinski||1651||Ozalj|1703||Graz|||
